library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;

entity bloque_6 is
end bloque_6 ;

architecture behavioral of bloque_6 is

begin


end behavioral;

